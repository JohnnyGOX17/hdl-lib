library ieee;
  use ieee.std_logic_1164.all;

entity cordic is
  generic (
    G_DATA_WIDTH : integer := 16
  );
  port (
    clk          : in  std_logic

  );
end entity cordic;

architecture rtl of cordic is

begin

end architecture rtl;
